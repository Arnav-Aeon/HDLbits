`timescale 1ns / 1ns
`include "2to1MUX.v"

module multiplex_gatelevel;

multiplex_gatelevel(z)

endmodule
